`timescale  1ns/1ns


module  vga_pic
(
    input   wire            vga_clk     ,   
    input   wire            sys_rst_n   ,   
    input   wire    [9:0]   pix_x       ,   
    input   wire    [9:0]   pix_y       ,   

    output  reg     [15:0]  pix_data        
);

parameter   CHAR_B_H=   10'd192 ,   
            CHAR_B_V=   10'd208 ;   

parameter   CHAR_W  =   10'd256 ,   
            CHAR_H  =   10'd64  ;   

parameter   BLACK   =   16'h0000,   
            WHITE   =   16'hFFFF,   
            GOLDEN  =   16'hFEC0;   


wire    [9:0]   char_x  ;   
wire    [9:0]   char_y  ;   

reg     [255:0] char    [63:0]  ;   

assign  char_x  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_x - CHAR_B_H) : 10'h3FF;
assign  char_y  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_y - CHAR_B_V) : 10'h3FF;


always@(posedge vga_clk)
    begin
        char[0]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[1]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[2]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[3]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[4]     <=  256'h00000000003C0000000000000000000000000000000070000000000000000000;
        char[5]     <=  256'h0000000E003E00000000000000000000000000000000F0000000000000000000;
        char[6]     <=  256'h000000FF001F00000000000000000000000000000001F0000000000000400000;
        char[7]     <=  256'h000007FF000F00000000000000000000000010000001F8000000000000E00000;
        char[8]     <=  256'h00007FFE000F000000000000000000000003FE000001F8000000000000F00000;
        char[9]     <=  256'h0000FE7E003F00000000000000000000000FFF800001F80000003E0000F00000;
        char[10]    <=  256'h0000E07C01F8000000000000000000000007FF81F801FC0000003F0000F00000;
        char[11]    <=  256'h0000E0F80380000000000000000000000003FF80FE00780000003F0001E00000;
        char[12]    <=  256'h0000E0F80380000000000000000000000001FF80FF00780000003F0001E00000;
        char[13]    <=  256'h0780E1F003FC000000000000000000000000FF80FF80780000003E0001E00000;
        char[14]    <=  256'h07C0FFF003FE0000000000020000000000003F007F80780000003E0001E00000;
        char[15]    <=  256'h07E0FFE001FE0000000000070000000000000E007F00780000003C0001FF0000;
        char[16]    <=  256'h07F3FFE0000E00000000000700000000000000007E00F80000003C0001FF0000;
        char[17]    <=  256'h07F9FFC0000E00000000000F0000000000003E00CC01F80000007C0003FE0000;
        char[18]    <=  256'h03F9FFC0001C03E00000000F8000000000003F010001F80000007E0003F80000;
        char[19]    <=  256'h03F9FF8000781FF80000001F8000000000007F038001F8000000FF0007F00000;
        char[20]    <=  256'h03F9FF8001F07FF80000001F878000000000FE078001F8000000FF000FE00000;
        char[21]    <=  256'h03FDFF0007C3FFF00000003FFFC000000001FC07C001F8000001FF003FE00000;
        char[22]    <=  256'h03FDFF000F9F8FF00001C03FFFC000000007F807F001F8000007FE003FC00000;
        char[23]    <=  256'h03FFFE001FFF8FE00001E07FFFC00000001FF807FC01F800000FFC0003C00000;
        char[24]    <=  256'h01FFF0007FFF8FC00003E07FFC000000067FF007FE01FC00001FF80003800000;
        char[25]    <=  256'h01FFC000FFEF9F800003E0FE000000000FFFF003FC01FE00007FF00007800000;
        char[26]    <=  256'h01FF8001FF8F9F000007E0FE000000000FFFF041F803FC0000FFE00007800000;
        char[27]    <=  256'h01FF8007FC1F9E00001FE0FE000000000FFFF180F00FFC000001E00007000000;
        char[28]    <=  256'h00FF8007F01F3C00003FE1FC00000000007FF601E01FF8000001E000071C0000;
        char[29]    <=  256'h00FF8007C01FFC00003FE1FC00000000001FFC03C0FFF8000001E0000F3E0000;
        char[30]    <=  256'h00030002001FF800003FC3FC00000000003FF807C3FFF8000001E7800FFE0000;
        char[31]    <=  256'h00070000001FF000007FC3F800000000003FF80F9FFFF0000001FF000FFE0000;
        char[32]    <=  256'h0007F000001FE000007F83F800000000007FF01FFFC3F0000001FE000FFE0000;
        char[33]    <=  256'h001FF000001FC000003F83F00000000000FFF01FFE03F0000001FC001FFE0000;
        char[34]    <=  256'h007FE000001F8000003F07F00000000000FFE03FF003F0000003F8001F3E0000;
        char[35]    <=  256'h007FC000001F8000001807F00000000001FFE03F8003F0000003F0001F3C0000;
        char[36]    <=  256'h00078600001F000000000FF80000000003FFC07E0003F0000003F0001E3C0000;
        char[37]    <=  256'h000F1E00001F000000000FFC0000000007FFC0180003F0000007E003843C0000;
        char[38]    <=  256'h003FFC00001F800000001FDE0000000007FFC0000003F000000FF001E03C0000;
        char[39]    <=  256'h007FF800001F800000003FDF8000000007C7C0000003F00000FFF000F83C0000;
        char[40]    <=  256'h00FFF000001F800000007F9FF00000000787C0000003F00007FFF0007F3C0000;
        char[41]    <=  256'h01FFE000001F80000000FF0FFE0000000707C0000003F0001FF1F8003FFC0000;
        char[42]    <=  256'h03FF8000001F80000001FE0FFFE000000003C0000003F0003F81F8001FFC0000;
        char[43]    <=  256'h07FF0000003F80000003FC07FFFE0000000300000003F0003E01FC000FFE0000;
        char[44]    <=  256'h07FC0000003F80000007F803FFFFE000000000000003F0001F83FC0007FFF000;
        char[45]    <=  256'h07F80000003F8000000FF001FFFFFF80000000000003F0000FFFFC0003FFFF80;
        char[46]    <=  256'h03E00000007F8000001FC0007FFFFFC0000000000003F00003FFFE0007FFFFF0;
        char[47]    <=  256'h0000000000FF8000007F80001FFFFFE0000000000003F000007FFE003FBFFFF8;
        char[48]    <=  256'h0000000001FF800000FE000007FFFFE0000000000003E000000FFC03FE0FFFF8;
        char[49]    <=  256'h0000000007FF800001F8000001FFFFF0000000000003E0000000F8FFC003FFF8;
        char[50]    <=  256'h000000007FFF000003E00000001FFFC0000000000003C0000000000000007FF8;
        char[51]    <=  256'h00000007FFFE0000070000000001FFC0000000000003C0000000000000000FF0;
        char[52]    <=  256'h0000000200F800000000000000000F8000000000000300000000000000000060;
        char[53]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[54]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[55]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[56]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[57]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[58]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[59]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[60]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[61]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[62]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[63]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
    end

always@(posedge vga_clk or negedge sys_rst_n)
    if(sys_rst_n == 1'b0)
        pix_data    <= BLACK;
    else    if((((pix_x >= (CHAR_B_H - 1'b1))
                && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
                && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                && (char[char_y][10'd255 - char_x] == 1'b1))
        pix_data    <=  GOLDEN;
    else
        pix_data    <=  BLACK;

endmodule
